//------------------------------------------------------
// Copyright 1992 Cascade Design Automation Corporation.
//------------------------------------------------------
module pd_wire(INN,INN);
  inout  INN;
endmodule
