//------------------------------------------------------
// Copyright 1992, 1993 Cascade Design Automation Corporation.
//------------------------------------------------------
module bufinv(IN0,Y);
  parameter N = 8;
  parameter DPFLAG = 0;
  parameter GROUP = "std";
  parameter
        d_IN0 = 0,
        d_Y = 1;
  input [(N - 1):0] IN0;
  output [(N - 1):0] Y;
  wire [(N - 1):0] IN0_temp;
  reg [(N - 1):0] Y_temp;
  assign #(d_IN0) IN0_temp = IN0;
  assign #(d_Y) Y = Y_temp;
  initial
    begin
    if((DPFLAG == 1))
      $display("(WARNING) The instance %m of type bufinv can't be implemented as a data-path cell");
    end
  always
    @(IN0_temp)
      Y_temp = ( ~ IN0_temp);
endmodule
